
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "seq_loop_interface.svh"
`include "seq_loop_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);




    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_top_kernel.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_top_kernel.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_top_kernel.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_103_1_fu_1199.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_103_1_fu_1199.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_103_1_fu_1199.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_2_VITIS_LOOP_110_3_fu_1235.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_2_VITIS_LOOP_110_3_fu_1235.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_2_VITIS_LOOP_110_3_fu_1235.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_5_fu_326.ap_start;
    assign module_intf_5.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_5_fu_326.ap_ready;
    assign module_intf_5.ap_done = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_5_fu_326.ap_done;
    assign module_intf_5.ap_continue = 1'b1;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_51_fu_364.ap_start;
    assign module_intf_6.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_51_fu_364.ap_ready;
    assign module_intf_6.ap_done = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_51_fu_364.ap_done;
    assign module_intf_6.ap_continue = 1'b1;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;
    nodf_module_intf module_intf_7(clock,reset);
    assign module_intf_7.ap_start = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_53_fu_402.ap_start;
    assign module_intf_7.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_53_fu_402.ap_ready;
    assign module_intf_7.ap_done = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_53_fu_402.ap_done;
    assign module_intf_7.ap_continue = 1'b1;
    assign module_intf_7.finish = finish;
    csv_file_dump mstatus_csv_dumper_7;
    nodf_module_monitor module_monitor_7;
    nodf_module_intf module_intf_8(clock,reset);
    assign module_intf_8.ap_start = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_55_fu_440.ap_start;
    assign module_intf_8.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_55_fu_440.ap_ready;
    assign module_intf_8.ap_done = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_55_fu_440.ap_done;
    assign module_intf_8.ap_continue = 1'b1;
    assign module_intf_8.finish = finish;
    csv_file_dump mstatus_csv_dumper_8;
    nodf_module_monitor module_monitor_8;
    nodf_module_intf module_intf_9(clock,reset);
    assign module_intf_9.ap_start = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_6_fu_478.ap_start;
    assign module_intf_9.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_6_fu_478.ap_ready;
    assign module_intf_9.ap_done = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_6_fu_478.ap_done;
    assign module_intf_9.ap_continue = 1'b1;
    assign module_intf_9.finish = finish;
    csv_file_dump mstatus_csv_dumper_9;
    nodf_module_monitor module_monitor_9;
    nodf_module_intf module_intf_10(clock,reset);
    assign module_intf_10.ap_start = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_62_fu_548.ap_start;
    assign module_intf_10.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_62_fu_548.ap_ready;
    assign module_intf_10.ap_done = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_62_fu_548.ap_done;
    assign module_intf_10.ap_continue = 1'b1;
    assign module_intf_10.finish = finish;
    csv_file_dump mstatus_csv_dumper_10;
    nodf_module_monitor module_monitor_10;
    nodf_module_intf module_intf_11(clock,reset);
    assign module_intf_11.ap_start = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_64_fu_618.ap_start;
    assign module_intf_11.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_64_fu_618.ap_ready;
    assign module_intf_11.ap_done = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_64_fu_618.ap_done;
    assign module_intf_11.ap_continue = 1'b1;
    assign module_intf_11.finish = finish;
    csv_file_dump mstatus_csv_dumper_11;
    nodf_module_monitor module_monitor_11;
    nodf_module_intf module_intf_12(clock,reset);
    assign module_intf_12.ap_start = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_66_fu_688.ap_start;
    assign module_intf_12.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_66_fu_688.ap_ready;
    assign module_intf_12.ap_done = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_66_fu_688.ap_done;
    assign module_intf_12.ap_continue = 1'b1;
    assign module_intf_12.finish = finish;
    csv_file_dump mstatus_csv_dumper_12;
    nodf_module_monitor module_monitor_12;
    nodf_module_intf module_intf_13(clock,reset);
    assign module_intf_13.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_139_7_VITIS_LOOP_140_8_fu_1438.ap_start;
    assign module_intf_13.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_139_7_VITIS_LOOP_140_8_fu_1438.ap_ready;
    assign module_intf_13.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_139_7_VITIS_LOOP_140_8_fu_1438.ap_done;
    assign module_intf_13.ap_continue = 1'b1;
    assign module_intf_13.finish = finish;
    csv_file_dump mstatus_csv_dumper_13;
    nodf_module_monitor module_monitor_13;
    nodf_module_intf module_intf_14(clock,reset);
    assign module_intf_14.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_10_fu_1522.ap_start;
    assign module_intf_14.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_10_fu_1522.ap_ready;
    assign module_intf_14.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_10_fu_1522.ap_done;
    assign module_intf_14.ap_continue = 1'b1;
    assign module_intf_14.finish = finish;
    csv_file_dump mstatus_csv_dumper_14;
    nodf_module_monitor module_monitor_14;
    nodf_module_intf module_intf_15(clock,reset);
    assign module_intf_15.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_107_fu_1561.ap_start;
    assign module_intf_15.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_107_fu_1561.ap_ready;
    assign module_intf_15.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_107_fu_1561.ap_done;
    assign module_intf_15.ap_continue = 1'b1;
    assign module_intf_15.finish = finish;
    csv_file_dump mstatus_csv_dumper_15;
    nodf_module_monitor module_monitor_15;
    nodf_module_intf module_intf_16(clock,reset);
    assign module_intf_16.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_108_fu_1600.ap_start;
    assign module_intf_16.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_108_fu_1600.ap_ready;
    assign module_intf_16.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_108_fu_1600.ap_done;
    assign module_intf_16.ap_continue = 1'b1;
    assign module_intf_16.finish = finish;
    csv_file_dump mstatus_csv_dumper_16;
    nodf_module_monitor module_monitor_16;
    nodf_module_intf module_intf_17(clock,reset);
    assign module_intf_17.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_109_fu_1639.ap_start;
    assign module_intf_17.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_109_fu_1639.ap_ready;
    assign module_intf_17.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_109_fu_1639.ap_done;
    assign module_intf_17.ap_continue = 1'b1;
    assign module_intf_17.finish = finish;
    csv_file_dump mstatus_csv_dumper_17;
    nodf_module_monitor module_monitor_17;
    nodf_module_intf module_intf_18(clock,reset);
    assign module_intf_18.ap_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_160_11_VITIS_LOOP_161_12_fu_1678.ap_start;
    assign module_intf_18.ap_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_160_11_VITIS_LOOP_161_12_fu_1678.ap_ready;
    assign module_intf_18.ap_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_160_11_VITIS_LOOP_161_12_fu_1678.ap_done;
    assign module_intf_18.ap_continue = 1'b1;
    assign module_intf_18.finish = finish;
    csv_file_dump mstatus_csv_dumper_18;
    nodf_module_monitor module_monitor_18;

    seq_loop_intf#(26) seq_loop_intf_1(clock,reset);
    assign seq_loop_intf_1.pre_loop_state0 = AESL_inst_top_kernel.ap_ST_fsm_state16;
    assign seq_loop_intf_1.pre_states_valid = 1'b1;
    assign seq_loop_intf_1.post_loop_state0 = AESL_inst_top_kernel.ap_ST_fsm_state20;
    assign seq_loop_intf_1.post_states_valid = 1'b1;
    assign seq_loop_intf_1.quit_loop_state0 = AESL_inst_top_kernel.ap_ST_fsm_state17;
    assign seq_loop_intf_1.quit_states_valid = 1'b1;
    assign seq_loop_intf_1.cur_state = AESL_inst_top_kernel.ap_CS_fsm;
    assign seq_loop_intf_1.iter_start_state = AESL_inst_top_kernel.ap_ST_fsm_state17;
    assign seq_loop_intf_1.iter_end_state0 = AESL_inst_top_kernel.ap_ST_fsm_state19;
    assign seq_loop_intf_1.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_1.one_state_loop = 1'b0;
    assign seq_loop_intf_1.one_state_block = 1'b0;
    assign seq_loop_intf_1.finish = finish;
    csv_file_dump seq_loop_csv_dumper_1;
    seq_loop_monitor #(26) seq_loop_monitor_1;
    seq_loop_intf#(5) seq_loop_intf_2(clock,reset);
    assign seq_loop_intf_2.pre_loop_state0 = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.ap_ST_fsm_state1;
    assign seq_loop_intf_2.pre_states_valid = 1'b1;
    assign seq_loop_intf_2.post_loop_state0 = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.ap_ST_fsm_state1;
    assign seq_loop_intf_2.post_states_valid = 1'b1;
    assign seq_loop_intf_2.quit_loop_state0 = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.ap_ST_fsm_state2;
    assign seq_loop_intf_2.quit_states_valid = 1'b1;
    assign seq_loop_intf_2.cur_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.ap_CS_fsm;
    assign seq_loop_intf_2.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.ap_ST_fsm_state2;
    assign seq_loop_intf_2.iter_end_state0 = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.ap_ST_fsm_state5;
    assign seq_loop_intf_2.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_2.one_state_loop = 1'b0;
    assign seq_loop_intf_2.one_state_block = 1'b0;
    assign seq_loop_intf_2.finish = finish;
    csv_file_dump seq_loop_csv_dumper_2;
    seq_loop_monitor #(5) seq_loop_monitor_2;
    upc_loop_intf#(1) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_103_1_fu_1199.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_103_1_fu_1199.ap_ST_fsm_state1;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_103_1_fu_1199.ap_ST_fsm_state1;
    assign upc_loop_intf_1.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_103_1_fu_1199.ap_ST_fsm_state1;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_103_1_fu_1199.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_103_1_fu_1199.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_1.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_103_1_fu_1199.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_1.iter_start_enable = 1'b1;
    assign upc_loop_intf_1.iter_end_enable = 1'b1;
    assign upc_loop_intf_1.quit_enable = 1'b1;
    assign upc_loop_intf_1.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_103_1_fu_1199.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_103_1_fu_1199.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_103_1_fu_1199.ap_done_int;
    assign upc_loop_intf_1.loop_continue = 1'b1;
    assign upc_loop_intf_1.quit_at_end = 1'b1;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(1) upc_loop_monitor_1;
    upc_loop_intf#(1) upc_loop_intf_2(clock,reset);
    assign upc_loop_intf_2.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_2_VITIS_LOOP_110_3_fu_1235.ap_CS_fsm;
    assign upc_loop_intf_2.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_2_VITIS_LOOP_110_3_fu_1235.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_2_VITIS_LOOP_110_3_fu_1235.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_2_VITIS_LOOP_110_3_fu_1235.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_2_VITIS_LOOP_110_3_fu_1235.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_2_VITIS_LOOP_110_3_fu_1235.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_2_VITIS_LOOP_110_3_fu_1235.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_2_VITIS_LOOP_110_3_fu_1235.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_2.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_2_VITIS_LOOP_110_3_fu_1235.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_2.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_2_VITIS_LOOP_110_3_fu_1235.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_2.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_2_VITIS_LOOP_110_3_fu_1235.ap_start;
    assign upc_loop_intf_2.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_2_VITIS_LOOP_110_3_fu_1235.ap_ready;
    assign upc_loop_intf_2.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_109_2_VITIS_LOOP_110_3_fu_1235.ap_done_int;
    assign upc_loop_intf_2.loop_continue = 1'b1;
    assign upc_loop_intf_2.quit_at_end = 1'b1;
    assign upc_loop_intf_2.finish = finish;
    csv_file_dump upc_loop_csv_dumper_2;
    upc_loop_monitor #(1) upc_loop_monitor_2;
    upc_loop_intf#(1) upc_loop_intf_3(clock,reset);
    assign upc_loop_intf_3.cur_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_5_fu_326.ap_CS_fsm;
    assign upc_loop_intf_3.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_5_fu_326.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_5_fu_326.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.quit_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_5_fu_326.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_5_fu_326.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_5_fu_326.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.quit_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_5_fu_326.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_5_fu_326.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_3.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_5_fu_326.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_3.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_5_fu_326.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_3.loop_start = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_5_fu_326.ap_start;
    assign upc_loop_intf_3.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_5_fu_326.ap_ready;
    assign upc_loop_intf_3.loop_done = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_5_fu_326.ap_done_int;
    assign upc_loop_intf_3.loop_continue = 1'b1;
    assign upc_loop_intf_3.quit_at_end = 1'b1;
    assign upc_loop_intf_3.finish = finish;
    csv_file_dump upc_loop_csv_dumper_3;
    upc_loop_monitor #(1) upc_loop_monitor_3;
    upc_loop_intf#(1) upc_loop_intf_4(clock,reset);
    assign upc_loop_intf_4.cur_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_51_fu_364.ap_CS_fsm;
    assign upc_loop_intf_4.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_51_fu_364.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_51_fu_364.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.quit_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_51_fu_364.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_51_fu_364.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_51_fu_364.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.quit_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_51_fu_364.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_51_fu_364.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_4.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_51_fu_364.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_4.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_51_fu_364.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_4.loop_start = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_51_fu_364.ap_start;
    assign upc_loop_intf_4.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_51_fu_364.ap_ready;
    assign upc_loop_intf_4.loop_done = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_51_fu_364.ap_done_int;
    assign upc_loop_intf_4.loop_continue = 1'b1;
    assign upc_loop_intf_4.quit_at_end = 1'b1;
    assign upc_loop_intf_4.finish = finish;
    csv_file_dump upc_loop_csv_dumper_4;
    upc_loop_monitor #(1) upc_loop_monitor_4;
    upc_loop_intf#(1) upc_loop_intf_5(clock,reset);
    assign upc_loop_intf_5.cur_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_53_fu_402.ap_CS_fsm;
    assign upc_loop_intf_5.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_53_fu_402.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_53_fu_402.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.quit_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_53_fu_402.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_53_fu_402.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_53_fu_402.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.quit_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_53_fu_402.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_53_fu_402.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_5.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_53_fu_402.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_5.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_53_fu_402.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_5.loop_start = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_53_fu_402.ap_start;
    assign upc_loop_intf_5.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_53_fu_402.ap_ready;
    assign upc_loop_intf_5.loop_done = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_53_fu_402.ap_done_int;
    assign upc_loop_intf_5.loop_continue = 1'b1;
    assign upc_loop_intf_5.quit_at_end = 1'b1;
    assign upc_loop_intf_5.finish = finish;
    csv_file_dump upc_loop_csv_dumper_5;
    upc_loop_monitor #(1) upc_loop_monitor_5;
    upc_loop_intf#(1) upc_loop_intf_6(clock,reset);
    assign upc_loop_intf_6.cur_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_55_fu_440.ap_CS_fsm;
    assign upc_loop_intf_6.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_55_fu_440.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_55_fu_440.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.quit_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_55_fu_440.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_55_fu_440.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_55_fu_440.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.quit_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_55_fu_440.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_55_fu_440.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_55_fu_440.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_6.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_55_fu_440.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_6.loop_start = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_55_fu_440.ap_start;
    assign upc_loop_intf_6.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_55_fu_440.ap_ready;
    assign upc_loop_intf_6.loop_done = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_121_55_fu_440.ap_done_int;
    assign upc_loop_intf_6.loop_continue = 1'b1;
    assign upc_loop_intf_6.quit_at_end = 1'b1;
    assign upc_loop_intf_6.finish = finish;
    csv_file_dump upc_loop_csv_dumper_6;
    upc_loop_monitor #(1) upc_loop_monitor_6;
    upc_loop_intf#(1) upc_loop_intf_7(clock,reset);
    assign upc_loop_intf_7.cur_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_6_fu_478.ap_CS_fsm;
    assign upc_loop_intf_7.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_6_fu_478.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_6_fu_478.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.quit_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_6_fu_478.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_6_fu_478.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_6_fu_478.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.quit_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_6_fu_478.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_6_fu_478.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_7.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_6_fu_478.ap_enable_reg_pp0_iter42;
    assign upc_loop_intf_7.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_6_fu_478.ap_enable_reg_pp0_iter42;
    assign upc_loop_intf_7.loop_start = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_6_fu_478.ap_start;
    assign upc_loop_intf_7.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_6_fu_478.ap_ready;
    assign upc_loop_intf_7.loop_done = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_6_fu_478.ap_done_int;
    assign upc_loop_intf_7.loop_continue = 1'b1;
    assign upc_loop_intf_7.quit_at_end = 1'b1;
    assign upc_loop_intf_7.finish = finish;
    csv_file_dump upc_loop_csv_dumper_7;
    upc_loop_monitor #(1) upc_loop_monitor_7;
    upc_loop_intf#(1) upc_loop_intf_8(clock,reset);
    assign upc_loop_intf_8.cur_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_62_fu_548.ap_CS_fsm;
    assign upc_loop_intf_8.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_62_fu_548.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_62_fu_548.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.quit_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_62_fu_548.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_62_fu_548.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_62_fu_548.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.quit_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_62_fu_548.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_62_fu_548.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_8.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_62_fu_548.ap_enable_reg_pp0_iter42;
    assign upc_loop_intf_8.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_62_fu_548.ap_enable_reg_pp0_iter42;
    assign upc_loop_intf_8.loop_start = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_62_fu_548.ap_start;
    assign upc_loop_intf_8.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_62_fu_548.ap_ready;
    assign upc_loop_intf_8.loop_done = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_62_fu_548.ap_done_int;
    assign upc_loop_intf_8.loop_continue = 1'b1;
    assign upc_loop_intf_8.quit_at_end = 1'b1;
    assign upc_loop_intf_8.finish = finish;
    csv_file_dump upc_loop_csv_dumper_8;
    upc_loop_monitor #(1) upc_loop_monitor_8;
    upc_loop_intf#(1) upc_loop_intf_9(clock,reset);
    assign upc_loop_intf_9.cur_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_64_fu_618.ap_CS_fsm;
    assign upc_loop_intf_9.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_64_fu_618.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_64_fu_618.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.quit_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_64_fu_618.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_64_fu_618.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_64_fu_618.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.quit_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_64_fu_618.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_64_fu_618.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_9.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_64_fu_618.ap_enable_reg_pp0_iter42;
    assign upc_loop_intf_9.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_64_fu_618.ap_enable_reg_pp0_iter42;
    assign upc_loop_intf_9.loop_start = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_64_fu_618.ap_start;
    assign upc_loop_intf_9.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_64_fu_618.ap_ready;
    assign upc_loop_intf_9.loop_done = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_64_fu_618.ap_done_int;
    assign upc_loop_intf_9.loop_continue = 1'b1;
    assign upc_loop_intf_9.quit_at_end = 1'b1;
    assign upc_loop_intf_9.finish = finish;
    csv_file_dump upc_loop_csv_dumper_9;
    upc_loop_monitor #(1) upc_loop_monitor_9;
    upc_loop_intf#(1) upc_loop_intf_10(clock,reset);
    assign upc_loop_intf_10.cur_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_66_fu_688.ap_CS_fsm;
    assign upc_loop_intf_10.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_66_fu_688.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_66_fu_688.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.quit_state = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_66_fu_688.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_66_fu_688.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_66_fu_688.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.quit_block = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_66_fu_688.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_66_fu_688.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_10.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_66_fu_688.ap_enable_reg_pp0_iter42;
    assign upc_loop_intf_10.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_66_fu_688.ap_enable_reg_pp0_iter42;
    assign upc_loop_intf_10.loop_start = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_66_fu_688.ap_start;
    assign upc_loop_intf_10.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_66_fu_688.ap_ready;
    assign upc_loop_intf_10.loop_done = AESL_inst_top_kernel.grp_top_kernel_Outline_VITIS_LOOP_117_4_fu_1306.grp_top_kernel_Pipeline_VITIS_LOOP_129_66_fu_688.ap_done_int;
    assign upc_loop_intf_10.loop_continue = 1'b1;
    assign upc_loop_intf_10.quit_at_end = 1'b1;
    assign upc_loop_intf_10.finish = finish;
    csv_file_dump upc_loop_csv_dumper_10;
    upc_loop_monitor #(1) upc_loop_monitor_10;
    upc_loop_intf#(1) upc_loop_intf_11(clock,reset);
    assign upc_loop_intf_11.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_139_7_VITIS_LOOP_140_8_fu_1438.ap_CS_fsm;
    assign upc_loop_intf_11.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_139_7_VITIS_LOOP_140_8_fu_1438.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_139_7_VITIS_LOOP_140_8_fu_1438.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_139_7_VITIS_LOOP_140_8_fu_1438.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_139_7_VITIS_LOOP_140_8_fu_1438.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_139_7_VITIS_LOOP_140_8_fu_1438.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_139_7_VITIS_LOOP_140_8_fu_1438.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_139_7_VITIS_LOOP_140_8_fu_1438.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_11.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_139_7_VITIS_LOOP_140_8_fu_1438.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_11.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_139_7_VITIS_LOOP_140_8_fu_1438.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_11.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_139_7_VITIS_LOOP_140_8_fu_1438.ap_start;
    assign upc_loop_intf_11.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_139_7_VITIS_LOOP_140_8_fu_1438.ap_ready;
    assign upc_loop_intf_11.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_139_7_VITIS_LOOP_140_8_fu_1438.ap_done_int;
    assign upc_loop_intf_11.loop_continue = 1'b1;
    assign upc_loop_intf_11.quit_at_end = 1'b1;
    assign upc_loop_intf_11.finish = finish;
    csv_file_dump upc_loop_csv_dumper_11;
    upc_loop_monitor #(1) upc_loop_monitor_11;
    upc_loop_intf#(2) upc_loop_intf_12(clock,reset);
    assign upc_loop_intf_12.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_10_fu_1522.ap_CS_fsm;
    assign upc_loop_intf_12.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_10_fu_1522.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_10_fu_1522.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_12.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_10_fu_1522.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_12.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_10_fu_1522.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_10_fu_1522.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_12.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_10_fu_1522.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_12.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_10_fu_1522.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_12.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_10_fu_1522.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_12.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_10_fu_1522.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_12.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_10_fu_1522.ap_start;
    assign upc_loop_intf_12.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_10_fu_1522.ap_ready;
    assign upc_loop_intf_12.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_10_fu_1522.ap_done_int;
    assign upc_loop_intf_12.loop_continue = 1'b1;
    assign upc_loop_intf_12.quit_at_end = 1'b1;
    assign upc_loop_intf_12.finish = finish;
    csv_file_dump upc_loop_csv_dumper_12;
    upc_loop_monitor #(2) upc_loop_monitor_12;
    upc_loop_intf#(2) upc_loop_intf_13(clock,reset);
    assign upc_loop_intf_13.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_107_fu_1561.ap_CS_fsm;
    assign upc_loop_intf_13.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_107_fu_1561.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_107_fu_1561.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_13.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_107_fu_1561.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_13.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_107_fu_1561.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_107_fu_1561.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_13.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_107_fu_1561.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_13.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_107_fu_1561.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_13.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_107_fu_1561.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_13.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_107_fu_1561.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_13.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_107_fu_1561.ap_start;
    assign upc_loop_intf_13.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_107_fu_1561.ap_ready;
    assign upc_loop_intf_13.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_107_fu_1561.ap_done_int;
    assign upc_loop_intf_13.loop_continue = 1'b1;
    assign upc_loop_intf_13.quit_at_end = 1'b1;
    assign upc_loop_intf_13.finish = finish;
    csv_file_dump upc_loop_csv_dumper_13;
    upc_loop_monitor #(2) upc_loop_monitor_13;
    upc_loop_intf#(2) upc_loop_intf_14(clock,reset);
    assign upc_loop_intf_14.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_108_fu_1600.ap_CS_fsm;
    assign upc_loop_intf_14.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_108_fu_1600.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_108_fu_1600.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_14.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_108_fu_1600.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_14.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_108_fu_1600.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_108_fu_1600.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_14.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_108_fu_1600.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_14.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_108_fu_1600.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_14.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_108_fu_1600.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_14.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_108_fu_1600.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_14.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_108_fu_1600.ap_start;
    assign upc_loop_intf_14.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_108_fu_1600.ap_ready;
    assign upc_loop_intf_14.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_108_fu_1600.ap_done_int;
    assign upc_loop_intf_14.loop_continue = 1'b1;
    assign upc_loop_intf_14.quit_at_end = 1'b1;
    assign upc_loop_intf_14.finish = finish;
    csv_file_dump upc_loop_csv_dumper_14;
    upc_loop_monitor #(2) upc_loop_monitor_14;
    upc_loop_intf#(2) upc_loop_intf_15(clock,reset);
    assign upc_loop_intf_15.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_109_fu_1639.ap_CS_fsm;
    assign upc_loop_intf_15.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_109_fu_1639.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_109_fu_1639.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_15.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_109_fu_1639.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_15.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_109_fu_1639.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_109_fu_1639.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_15.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_109_fu_1639.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_15.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_109_fu_1639.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_15.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_109_fu_1639.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_15.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_109_fu_1639.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_15.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_109_fu_1639.ap_start;
    assign upc_loop_intf_15.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_109_fu_1639.ap_ready;
    assign upc_loop_intf_15.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_152_109_fu_1639.ap_done_int;
    assign upc_loop_intf_15.loop_continue = 1'b1;
    assign upc_loop_intf_15.quit_at_end = 1'b1;
    assign upc_loop_intf_15.finish = finish;
    csv_file_dump upc_loop_csv_dumper_15;
    upc_loop_monitor #(2) upc_loop_monitor_15;
    upc_loop_intf#(1) upc_loop_intf_16(clock,reset);
    assign upc_loop_intf_16.cur_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_160_11_VITIS_LOOP_161_12_fu_1678.ap_CS_fsm;
    assign upc_loop_intf_16.iter_start_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_160_11_VITIS_LOOP_161_12_fu_1678.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.iter_end_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_160_11_VITIS_LOOP_161_12_fu_1678.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.quit_state = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_160_11_VITIS_LOOP_161_12_fu_1678.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.iter_start_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_160_11_VITIS_LOOP_161_12_fu_1678.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.iter_end_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_160_11_VITIS_LOOP_161_12_fu_1678.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.quit_block = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_160_11_VITIS_LOOP_161_12_fu_1678.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.iter_start_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_160_11_VITIS_LOOP_161_12_fu_1678.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_16.iter_end_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_160_11_VITIS_LOOP_161_12_fu_1678.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_16.quit_enable = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_160_11_VITIS_LOOP_161_12_fu_1678.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_16.loop_start = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_160_11_VITIS_LOOP_161_12_fu_1678.ap_start;
    assign upc_loop_intf_16.loop_ready = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_160_11_VITIS_LOOP_161_12_fu_1678.ap_ready;
    assign upc_loop_intf_16.loop_done = AESL_inst_top_kernel.grp_top_kernel_Pipeline_VITIS_LOOP_160_11_VITIS_LOOP_161_12_fu_1678.ap_done_int;
    assign upc_loop_intf_16.loop_continue = 1'b1;
    assign upc_loop_intf_16.quit_at_end = 1'b1;
    assign upc_loop_intf_16.finish = finish;
    csv_file_dump upc_loop_csv_dumper_16;
    upc_loop_monitor #(1) upc_loop_monitor_16;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;



    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);
    mstatus_csv_dumper_7 = new("./module_status7.csv");
    module_monitor_7 = new(module_intf_7,mstatus_csv_dumper_7);
    mstatus_csv_dumper_8 = new("./module_status8.csv");
    module_monitor_8 = new(module_intf_8,mstatus_csv_dumper_8);
    mstatus_csv_dumper_9 = new("./module_status9.csv");
    module_monitor_9 = new(module_intf_9,mstatus_csv_dumper_9);
    mstatus_csv_dumper_10 = new("./module_status10.csv");
    module_monitor_10 = new(module_intf_10,mstatus_csv_dumper_10);
    mstatus_csv_dumper_11 = new("./module_status11.csv");
    module_monitor_11 = new(module_intf_11,mstatus_csv_dumper_11);
    mstatus_csv_dumper_12 = new("./module_status12.csv");
    module_monitor_12 = new(module_intf_12,mstatus_csv_dumper_12);
    mstatus_csv_dumper_13 = new("./module_status13.csv");
    module_monitor_13 = new(module_intf_13,mstatus_csv_dumper_13);
    mstatus_csv_dumper_14 = new("./module_status14.csv");
    module_monitor_14 = new(module_intf_14,mstatus_csv_dumper_14);
    mstatus_csv_dumper_15 = new("./module_status15.csv");
    module_monitor_15 = new(module_intf_15,mstatus_csv_dumper_15);
    mstatus_csv_dumper_16 = new("./module_status16.csv");
    module_monitor_16 = new(module_intf_16,mstatus_csv_dumper_16);
    mstatus_csv_dumper_17 = new("./module_status17.csv");
    module_monitor_17 = new(module_intf_17,mstatus_csv_dumper_17);
    mstatus_csv_dumper_18 = new("./module_status18.csv");
    module_monitor_18 = new(module_intf_18,mstatus_csv_dumper_18);



    seq_loop_csv_dumper_1 = new("./seq_loop_status1.csv");
    seq_loop_monitor_1 = new(seq_loop_intf_1,seq_loop_csv_dumper_1);
    seq_loop_csv_dumper_2 = new("./seq_loop_status2.csv");
    seq_loop_monitor_2 = new(seq_loop_intf_2,seq_loop_csv_dumper_2);

    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);
    upc_loop_csv_dumper_2 = new("./upc_loop_status2.csv");
    upc_loop_monitor_2 = new(upc_loop_intf_2,upc_loop_csv_dumper_2);
    upc_loop_csv_dumper_3 = new("./upc_loop_status3.csv");
    upc_loop_monitor_3 = new(upc_loop_intf_3,upc_loop_csv_dumper_3);
    upc_loop_csv_dumper_4 = new("./upc_loop_status4.csv");
    upc_loop_monitor_4 = new(upc_loop_intf_4,upc_loop_csv_dumper_4);
    upc_loop_csv_dumper_5 = new("./upc_loop_status5.csv");
    upc_loop_monitor_5 = new(upc_loop_intf_5,upc_loop_csv_dumper_5);
    upc_loop_csv_dumper_6 = new("./upc_loop_status6.csv");
    upc_loop_monitor_6 = new(upc_loop_intf_6,upc_loop_csv_dumper_6);
    upc_loop_csv_dumper_7 = new("./upc_loop_status7.csv");
    upc_loop_monitor_7 = new(upc_loop_intf_7,upc_loop_csv_dumper_7);
    upc_loop_csv_dumper_8 = new("./upc_loop_status8.csv");
    upc_loop_monitor_8 = new(upc_loop_intf_8,upc_loop_csv_dumper_8);
    upc_loop_csv_dumper_9 = new("./upc_loop_status9.csv");
    upc_loop_monitor_9 = new(upc_loop_intf_9,upc_loop_csv_dumper_9);
    upc_loop_csv_dumper_10 = new("./upc_loop_status10.csv");
    upc_loop_monitor_10 = new(upc_loop_intf_10,upc_loop_csv_dumper_10);
    upc_loop_csv_dumper_11 = new("./upc_loop_status11.csv");
    upc_loop_monitor_11 = new(upc_loop_intf_11,upc_loop_csv_dumper_11);
    upc_loop_csv_dumper_12 = new("./upc_loop_status12.csv");
    upc_loop_monitor_12 = new(upc_loop_intf_12,upc_loop_csv_dumper_12);
    upc_loop_csv_dumper_13 = new("./upc_loop_status13.csv");
    upc_loop_monitor_13 = new(upc_loop_intf_13,upc_loop_csv_dumper_13);
    upc_loop_csv_dumper_14 = new("./upc_loop_status14.csv");
    upc_loop_monitor_14 = new(upc_loop_intf_14,upc_loop_csv_dumper_14);
    upc_loop_csv_dumper_15 = new("./upc_loop_status15.csv");
    upc_loop_monitor_15 = new(upc_loop_intf_15,upc_loop_csv_dumper_15);
    upc_loop_csv_dumper_16 = new("./upc_loop_status16.csv");
    upc_loop_monitor_16 = new(upc_loop_intf_16,upc_loop_csv_dumper_16);

    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(module_monitor_7);
    sample_manager_inst.add_one_monitor(module_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_9);
    sample_manager_inst.add_one_monitor(module_monitor_10);
    sample_manager_inst.add_one_monitor(module_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_14);
    sample_manager_inst.add_one_monitor(module_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_16);
    sample_manager_inst.add_one_monitor(module_monitor_17);
    sample_manager_inst.add_one_monitor(module_monitor_18);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_1);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_2);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_2);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_3);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_4);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_5);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_6);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_7);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_8);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_9);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_10);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_11);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_12);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_13);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_14);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_15);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_16);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1) begin
                @(negedge clock);
                break;
            end
            else
                @(posedge clock);
        end
    endtask


endmodule
